A Berkeley SPICE3 compatible circuit  
*  
* This circuit contains only Berkeley SPICE3 components.  
*  
* The circuit is an AC coupled transistor amplifier with  
* a sinewave input at node "1", a gain of approximately -3.9,  
* and output on node "coll".  
*  
.tran 1e-5 2e-3  
*  
vcc vcc 0 12.0  
vin 1 0 0.0 ac 1.0 sin(0 1 1k)  
ccouple 1 base 10uF  
rbias1 vcc base 100k 
rbias2 base 0 24k  
q1 coll base emit generic
rcollector vcc coll 3.9k  
remitter emit 0 1k
*
.probe v(emit) v(vcc) v(1) v(base) v(coll) vcc#branch vin#branch
.model generic npn  
*    
.end